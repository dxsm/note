//------------------------------------------------------------------------
// File Name   : comb_shape.v
// Author      : victor dong (dxs_uestc@163.com)
// Version     : V0.1 
//------------------------------------------------------------------------
// Description :
//     
//------------------------------------------------------------------------
// Revision History:
// *Version* | *Modifier* | *Modified Date* | *Description*
//   V0.1    |   Victor   |   2019-10-20    | Fisrt Created.
//------------------------------------------------------------------------

module comb_shape(
  input               clk_a                   ,
  input               clk_b                   ,
  input               rst_a_n                 ,
  input               rst_b_n                 ,
  input               chip_head_in            ,

  //cell0 0~19 pool
  input               cell0_pool0_vld_in      ,
  input       [3:0]   cell0_pool0_chnum_in    ,
  input       [15:0]  cell0_pool0_data_in     ,
  input               cell0_pool0_10ms_timer  ,
  input               cell0_pool1_vld_in      ,
  input       [3:0]   cell0_pool1_chnum_in    ,
  input       [15:0]  cell0_pool1_data_in     ,
  input               cell0_pool1_10ms_timer  ,
  input               cell0_pool2_vld_in      ,
  input       [3:0]   cell0_pool2_chnum_in    ,
  input       [15:0]  cell0_pool2_data_in     ,
  input               cell0_pool2_10ms_timer  ,
  input               cell0_pool3_vld_in      ,
  input       [3:0]   cell0_pool3_chnum_in    ,
  input       [15:0]  cell0_pool3_data_in     ,
  input               cell0_pool3_10ms_timer  ,
  input               cell0_pool4_vld_in      ,
  input       [3:0]   cell0_pool4_chnum_in    ,
  input       [15:0]  cell0_pool4_data_in     ,
  input               cell0_pool4_10ms_timer  ,
  input               cell0_pool5_vld_in      ,
  input       [3:0]   cell0_pool5_chnum_in    ,
  input       [15:0]  cell0_pool5_data_in     ,
  input               cell0_pool5_10ms_timer  ,
  input               cell0_pool6_vld_in      ,
  input       [3:0]   cell0_pool6_chnum_in    ,
  input       [15:0]  cell0_pool6_data_in     ,
  input               cell0_pool6_10ms_timer  ,
  input               cell0_pool7_vld_in      ,
  input       [3:0]   cell0_pool7_chnum_in    ,
  input       [15:0]  cell0_pool0_data_in     ,
  input               cell0_pool0_10ms_timer  ,
  input               cell0_pool8_vld_in      ,
  input       [3:0]   cell0_pool8_chnum_in    ,
  input       [15:0]  cell0_pool8_data_in     ,
  input               cell0_pool8_10ms_timer  ,
  input               cell0_pool9_vld_in      ,
  input       [3:0]   cell0_pool9_chnum_in    ,
  input       [15:0]  cell0_pool9_data_in     ,
  input               cell0_pool9_10ms_timer  ,
  input               cell0_pool10_vld_in     ,
  input       [3:0]   cell0_pool10_chnum_in   ,
  input       [15:0]  cell0_pool10_data_in    ,
  input               cell0_pool10_10ms_timer ,
  input               cell0_pool11_vld_in     ,
  input       [3:0]   cell0_pool11_chnum_in   ,
  input       [15:0]  cell0_pool11_data_in    ,
  input               cell0_pool11_10ms_timer ,
  input               cell0_pool12_vld_in     ,
  input       [3:0]   cell0_pool12_chnum_in   ,
  input       [15:0]  cell0_pool12_data_in    ,
  input               cell0_pool12_10ms_timer ,
  input               cell0_pool13_vld_in     ,
  input       [3:0]   cell0_pool13_chnum_in   ,
  input       [15:0]  cell0_pool13_data_in    ,
  input               cell0_pool13_10ms_timer ,
  input               cell0_pool14_vld_in     ,
  input       [3:0]   cell0_pool14_chnum_in   ,
  input       [15:0]  cell0_pool14_data_in    ,
  input               cell0_pool14_10ms_timer ,
  input               cell0_pool15_vld_in     ,
  input       [3:0]   cell0_pool15_chnum_in   ,
  input       [15:0]  cell0_pool15_data_in    ,
  input               cell0_pool15_10ms_timer ,
  input               cell0_pool16_vld_in     ,
  input       [3:0]   cell0_pool16_chnum_in   ,
  input       [15:0]  cell0_pool16_data_in    ,
  input               cell0_pool16_10ms_timer ,
  input               cell0_pool17_vld_in     ,
  input       [3:0]   cell0_pool17_chnum_in   ,
  input       [15:0]  cell0_pool17_data_in    ,
  input               cell0_pool17_10ms_timer ,
  input               cell0_pool18_vld_in     ,
  input       [3:0]   cell0_pool18_chnum_in   ,
  input       [15:0]  cell0_pool18_data_in    ,
  input               cell0_pool18_10ms_timer ,
  input               cell0_pool19_vld_in     ,
  input       [3:0]   cell0_pool19_chnum_in   ,
  input       [15:0]  cell0_pool19_data_in    ,
  input               cell0_pool19_10ms_timer ,

  //cell1 0~19 pool
  input               cell1_pool0_vld_in      ,
  input       [3:0]   cell1_pool0_chnum_in    ,
  input       [15:0]  cell1_pool0_data_in     ,
  input               cell1_pool0_10ms_timer  ,
  input               cell1_pool1_vld_in      ,
  input       [3:0]   cell1_pool1_chnum_in    ,
  input       [15:0]  cell1_pool1_data_in     ,
  input               cell1_pool1_10ms_timer  ,
  input               cell1_pool2_vld_in      ,
  input       [3:0]   cell1_pool2_chnum_in    ,
  input       [15:0]  cell1_pool2_data_in     ,
  input               cell1_pool2_10ms_timer  ,
  input               cell1_pool3_vld_in      ,
  input       [3:0]   cell1_pool3_chnum_in    ,
  input       [15:0]  cell1_pool3_data_in     ,
  input               cell1_pool3_10ms_timer  ,
  input               cell1_pool4_vld_in      ,
  input       [3:0]   cell1_pool4_chnum_in    ,
  input       [15:0]  cell1_pool4_data_in     ,
  input               cell1_pool4_10ms_timer  ,
  input               cell1_pool5_vld_in      ,
  input       [3:0]   cell1_pool5_chnum_in    ,
  input       [15:0]  cell1_pool5_data_in     ,
  input               cell1_pool5_10ms_timer  ,
  input               cell1_pool6_vld_in      ,
  input       [3:0]   cell1_pool6_chnum_in    ,
  input       [15:0]  cell1_pool6_data_in     ,
  input               cell1_pool6_10ms_timer  ,
  input               cell1_pool7_vld_in      ,
  input       [3:0]   cell1_pool7_chnum_in    ,
  input       [15:0]  cell1_pool0_data_in     ,
  input               cell1_pool0_10ms_timer  ,
  input               cell1_pool8_vld_in      ,
  input       [3:0]   cell1_pool8_chnum_in    ,
  input       [15:0]  cell1_pool8_data_in     ,
  input               cell1_pool8_10ms_timer  ,
  input               cell1_pool9_vld_in      ,
  input       [3:0]   cell1_pool9_chnum_in    ,
  input       [15:0]  cell1_pool9_data_in     ,
  input               cell1_pool9_10ms_timer  ,
  input               cell1_pool10_vld_in     ,
  input       [3:0]   cell1_pool10_chnum_in   ,
  input       [15:0]  cell1_pool10_data_in    ,
  input               cell1_pool10_10ms_timer ,
  input               cell1_pool11_vld_in     ,
  input       [3:0]   cell1_pool11_chnum_in   ,
  input       [15:0]  cell1_pool11_data_in    ,
  input               cell1_pool11_10ms_timer ,
  input               cell1_pool12_vld_in     ,
  input       [3:0]   cell1_pool12_chnum_in   ,
  input       [15:0]  cell1_pool12_data_in    ,
  input               cell1_pool12_10ms_timer ,
  input               cell1_pool13_vld_in     ,
  input       [3:0]   cell1_pool13_chnum_in   ,
  input       [15:0]  cell1_pool13_data_in    ,
  input               cell1_pool13_10ms_timer ,
  input               cell1_pool14_vld_in     ,
  input       [3:0]   cell1_pool14_chnum_in   ,
  input       [15:0]  cell1_pool14_data_in    ,
  input               cell1_pool14_10ms_timer ,
  input               cell1_pool15_vld_in     ,
  input       [3:0]   cell1_pool15_chnum_in   ,
  input       [15:0]  cell1_pool15_data_in    ,
  input               cell1_pool15_10ms_timer ,
  input               cell1_pool16_vld_in     ,
  input       [3:0]   cell1_pool16_chnum_in   ,
  input       [15:0]  cell1_pool16_data_in    ,
  input               cell1_pool16_10ms_timer ,
  input               cell1_pool17_vld_in     ,
  input       [3:0]   cell1_pool17_chnum_in   ,
  input       [15:0]  cell1_pool17_data_in    ,
  input               cell1_pool17_10ms_timer ,
  input               cell1_pool18_vld_in     ,
  input       [3:0]   cell1_pool18_chnum_in   ,
  input       [15:0]  cell1_pool18_data_in    ,
  input               cell1_pool18_10ms_timer ,
  input               cell1_pool19_vld_in     ,
  input       [3:0]   cell1_pool19_chnum_in   ,
  input       [15:0]  cell1_pool19_data_in    ,
  input               cell1_pool19_10ms_timer ,

  //shape out 0~7 pool
  output wire         chip_head_out           ,
  output wire         shape_pool0_vld_out     ,
  output wire [8:0]   shape_pool0_chnum_out   ,
  output wire [15:0]  shape_pool0_data_out    ,
  output wire         shape_pool1_vld_out     ,
  output wire [8:0]   shape_pool1_chnum_out   ,
  output wire [15:0]  shape_pool1_data_out    ,
  output wire         shape_pool2_vld_out     ,
  output wire [8:0]   shape_pool2_chnum_out   ,
  output wire [15:0]  shape_pool2_data_out    ,
  output wire         shape_pool3_vld_out     ,
  output wire [8:0]   shape_pool3_chnum_out   ,
  output wire [15:0]  shape_pool3_data_out    ,
  output wire         shape_pool4_vld_out     ,
  output wire [8:0]   shape_pool4_chnum_out   ,
  output wire [15:0]  shape_pool4_data_out    ,
  output wire         shape_pool5_vld_out     ,
  output wire [8:0]   shape_pool5_chnum_out   ,
  output wire [15:0]  shape_pool5_data_out    ,
  output wire         shape_pool6_vld_out     ,
  output wire [8:0]   shape_pool6_chnum_out   ,
  output wire [15:0]  shape_pool6_data_out    ,
  output wire         shape_pool7_vld_out     ,
  output wire [8:0]   shape_pool7_chnum_out   ,
  output wire [15:0]  shape_pool7_data_out     
);

//==============================================
// Definition of regs and wires
//==============================================

//**********************************************
// Function
//**********************************************

endmodule
